
`timescale 1ns/1ps

`include "define.vh"

module vote(
    // output 
    output bit [1:0]    res,

    // input
    input  bit [1:0]    label_nn1,
    input  bit [1:0]    label_nn2,
    input  bit [1:0]    label_nn3,
    input  bit [1:0]    label_nn4, // new
    input  bit [1:0]    label_nn5  // new

);


    // --------------------------------------------------------------
    // Implement your design from here









endmodule
