    Mac OS X            	   2   �      �                                      ATTR       �   �   R                  �   R  com.dropbox.attributes   x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%��LǪ��}�L ����Vnk�T[[ �p�