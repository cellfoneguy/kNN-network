
`define  NUM_BIT        8
